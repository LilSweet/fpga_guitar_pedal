// constants_pack.sv
package constants_pack;
	localparam logic [31:0] PI_Q824 = 32'h03243F6A; // 52690912 in Q(8,24)
	localparam logic [31:0] GAIN_FACTOR_Q824 = 32'h28000000;
	// Add more constants, types, or functions as needed
endpackage

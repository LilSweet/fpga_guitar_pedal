`ifndef DEV_DEF
`define DEV_DEF

`define VENDOR_NAME "XILINX"
`define DEVICE_NAME "A7"

//`define LATTICE
//`define LCMXO3D
////`define LCMXO3LF
////`define MAX10

`endif